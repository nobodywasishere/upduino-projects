library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity text_buffer is
	port(
        clk : in std_logic;
        row : in unsigned(5 downto 0);
        col : in unsigned(5 downto 0);
        char : out unsigned(7 downto 0)
	);
end text_buffer;

architecture synth of text_buffer is

    signal addr : unsigned (11 downto 0) := (others => '0');

begin

    addr <= row & col;

    process (clk) begin
        if (rising_edge(clk)) then
            case addr is

                -- First row
                when "000000000000" => char <= "01000001";
                when "000000000001" => char <= "01000010";
                when "000000000010" => char <= "01000011";
                when "000000000011" => char <= "01000100";
                when "000000000100" => char <= "01000101";
                when "000000000101" => char <= "01000110";
                when "000000000110" => char <= "01000111";
                when "000000000111" => char <= "01001000";
                when "000000001000" => char <= "01001001";
                when "000000001001" => char <= "01001010";
                when "000000001010" => char <= "01001011";
                when "000000001011" => char <= "01001100";
                when "000000001100" => char <= "01001101";
                when "000000001101" => char <= "01001110";
                when "000000001110" => char <= "01001111";
                when "000000001111" => char <= "01010000";
                when "000000010000" => char <= "01010001";
                when "000000010001" => char <= "01010010";
                when "000000010010" => char <= "01010011";
                when "000000010011" => char <= "01010100";
                when "000000010100" => char <= "01010101";
                when "000000010101" => char <= "01010110";
                when "000000010110" => char <= "01010111";
                when "000000010111" => char <= "01011000";
                when "000000011000" => char <= "01011001";
                when "000000011001" => char <= "01011010";
                when "000000011010" => char <= "01011011";
                when "000000011011" => char <= "01011100";
                when "000000011100" => char <= "01011101";
                when "000000011101" => char <= "01011110";
                when "000000011110" => char <= "01011111";
                when "000000011111" => char <= "01011111";
                when "000000100000" => char <= "00000000";
                when "000000100001" => char <= "00000000";
                when "000000100010" => char <= "00000000";
                when "000000100011" => char <= "00000000";
                when "000000100100" => char <= "00000000";
                when "000000100101" => char <= "00000000";
                when "000000100110" => char <= "00000000";
                when "000000100111" => char <= "00000000";
                when "000000101000" => char <= "00000000";

                -- 1st column
                when "000001000000" => char <= "01000010";
                when "000010000000" => char <= "01000011";
                when "000011000000" => char <= "01000100";
                when "000100000000" => char <= "01000101";
                when "000101000000" => char <= "01000110";
                when "000110000000" => char <= "01000111";
                when "000111000000" => char <= "01001000";
                when "001000000000" => char <= "01001001";
                when "001001000000" => char <= "01001010";
                when "001010000000" => char <= "01001011";
                when "001011000000" => char <= "01001100";
                when "001100000000" => char <= "01001101";
                when "001101000000" => char <= "01001110";
                when "001110000000" => char <= "01001111";
                when "001111000000" => char <= "01010000";
                when "010000000000" => char <= "01010001";
                when "010001000000" => char <= "01010010";
                when "010010000000" => char <= "01010011";
                when "010011000000" => char <= "01010100";
                when "010100000000" => char <= "01010101";
                when "010101000000" => char <= "01010110";
                when "010110000000" => char <= "01010111";
                when "010111000000" => char <= "01011000";
                when "011000000000" => char <= "01011001";
                when "011001000000" => char <= "01011010";
                when "011010000000" => char <= "01011011";
                when "011011000000" => char <= "01011100";
                when "011100000000" => char <= "01011101";
                when "011101000000" => char <= "01011110";
                when "011110000000" => char <= "01011111";
                when "011111000000" => char <= "01011111";

                when         others => char <= "00000000";
            end case;
        end if;
    end process;

end;
