
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity text_rom is
	port(
        clk : in std_logic;
        row : in unsigned(5 downto 0);
        col : in unsigned(5 downto 0);
        char : out unsigned(7 downto 0)
	);
end text_rom;

architecture synth of text_rom is

    signal addr : unsigned (11 downto 0) := (others => '0');

begin

    addr <= row & col;

    process (clk) begin
        if (rising_edge(clk)) then
            case addr is
                when "000000000001" => char <= "00100000";	--  
                when "000000000010" => char <= "00100000";	--  
                when "000000000011" => char <= "00100000";	--  
                when "000000000100" => char <= "01000000";	-- @
                when "000000000101" => char <= "01000000";	-- @
                when "000000000110" => char <= "01000000";	-- @
                when "000000000111" => char <= "00100000";	--  
                when "000000001000" => char <= "00100000";	--  
                when "000000001001" => char <= "00100000";	--  
                when "000000001010" => char <= "00100000";	--  
                when "000000001011" => char <= "00100000";	--  
                when "000000001100" => char <= "00100000";	--  
                when "000000001101" => char <= "01000000";	-- @
                when "000000001110" => char <= "01000000";	-- @
                when "000000001111" => char <= "01000000";	-- @

                when "000001000001" => char <= "00100000";	--  
                when "000001000010" => char <= "01000000";	-- @
                when "000001000011" => char <= "01000000";	-- @
                when "000001000100" => char <= "01000000";	-- @
                when "000001000101" => char <= "01000000";	-- @
                when "000001000110" => char <= "01000000";	-- @
                when "000001000111" => char <= "01000000";	-- @
                when "000001001000" => char <= "01000000";	-- @
                when "000001001001" => char <= "00100000";	--  
                when "000001001010" => char <= "00100000";	--  
                when "000001001011" => char <= "01000000";	-- @
                when "000001001100" => char <= "01000000";	-- @
                when "000001001101" => char <= "01000000";	-- @
                when "000001001110" => char <= "01000000";	-- @
                when "000001001111" => char <= "01000000";	-- @
                when "000001010000" => char <= "01000000";	-- @
                when "000001010001" => char <= "01000000";	-- @

                when "000010000001" => char <= "01000000";	-- @
                when "000010000010" => char <= "01000000";	-- @
                when "000010000011" => char <= "01000000";	-- @
                when "000010000100" => char <= "01000000";	-- @
                when "000010000101" => char <= "01000000";	-- @
                when "000010000110" => char <= "01000000";	-- @
                when "000010000111" => char <= "01000000";	-- @
                when "000010001000" => char <= "01000000";	-- @
                when "000010001001" => char <= "01000000";	-- @
                when "000010001010" => char <= "01000000";	-- @
                when "000010001011" => char <= "01000000";	-- @
                when "000010001100" => char <= "01000000";	-- @
                when "000010001101" => char <= "01000000";	-- @
                when "000010001110" => char <= "01000000";	-- @
                when "000010001111" => char <= "01000000";	-- @
                when "000010010000" => char <= "01000000";	-- @
                when "000010010001" => char <= "01000000";	-- @
                when "000010010010" => char <= "01000000";	-- @

                when "000011000001" => char <= "01000000";	-- @
                when "000011000010" => char <= "01000000";	-- @
                when "000011000011" => char <= "01000000";	-- @
                when "000011000100" => char <= "01000000";	-- @
                when "000011000101" => char <= "01000000";	-- @
                when "000011000110" => char <= "01000000";	-- @
                when "000011000111" => char <= "01000000";	-- @
                when "000011001000" => char <= "01000000";	-- @
                when "000011001001" => char <= "01000000";	-- @
                when "000011001010" => char <= "01000000";	-- @
                when "000011001011" => char <= "01000000";	-- @
                when "000011001100" => char <= "01000000";	-- @
                when "000011001101" => char <= "01000000";	-- @
                when "000011001110" => char <= "01000000";	-- @
                when "000011001111" => char <= "01000000";	-- @
                when "000011010000" => char <= "01000000";	-- @
                when "000011010001" => char <= "01000000";	-- @
                when "000011010010" => char <= "01000000";	-- @

                when "000100000001" => char <= "01000000";	-- @
                when "000100000010" => char <= "01000000";	-- @
                when "000100000011" => char <= "01000000";	-- @
                when "000100000100" => char <= "01000000";	-- @
                when "000100000101" => char <= "01000000";	-- @
                when "000100000110" => char <= "01000000";	-- @
                when "000100000111" => char <= "01000000";	-- @
                when "000100001000" => char <= "01000000";	-- @
                when "000100001001" => char <= "01000000";	-- @
                when "000100001010" => char <= "01000000";	-- @
                when "000100001011" => char <= "01000000";	-- @
                when "000100001100" => char <= "01000000";	-- @
                when "000100001101" => char <= "01000000";	-- @
                when "000100001110" => char <= "01000000";	-- @
                when "000100001111" => char <= "01000000";	-- @
                when "000100010000" => char <= "01000000";	-- @
                when "000100010001" => char <= "01000000";	-- @
                when "000100010010" => char <= "01000000";	-- @

                when "000101000001" => char <= "00100000";	--  
                when "000101000010" => char <= "01000000";	-- @
                when "000101000011" => char <= "01000000";	-- @
                when "000101000100" => char <= "01000000";	-- @
                when "000101000101" => char <= "01000000";	-- @
                when "000101000110" => char <= "01000000";	-- @
                when "000101000111" => char <= "01000000";	-- @
                when "000101001000" => char <= "01000000";	-- @
                when "000101001001" => char <= "01000000";	-- @
                when "000101001010" => char <= "01000000";	-- @
                when "000101001011" => char <= "01000000";	-- @
                when "000101001100" => char <= "01000000";	-- @
                when "000101001101" => char <= "01000000";	-- @
                when "000101001110" => char <= "01000000";	-- @
                when "000101001111" => char <= "01000000";	-- @
                when "000101010000" => char <= "01000000";	-- @
                when "000101010001" => char <= "01000000";	-- @

                when "000110000001" => char <= "00100000";	--  
                when "000110000010" => char <= "00100000";	--  
                when "000110000011" => char <= "00100000";	--  
                when "000110000100" => char <= "01000000";	-- @
                when "000110000101" => char <= "01000000";	-- @
                when "000110000110" => char <= "01000000";	-- @
                when "000110000111" => char <= "01000000";	-- @
                when "000110001000" => char <= "01000000";	-- @
                when "000110001001" => char <= "01000000";	-- @
                when "000110001010" => char <= "01000000";	-- @
                when "000110001011" => char <= "01000000";	-- @
                when "000110001100" => char <= "01000000";	-- @
                when "000110001101" => char <= "01000000";	-- @
                when "000110001110" => char <= "01000000";	-- @
                when "000110001111" => char <= "01000000";	-- @

                when "000111000001" => char <= "00100000";	--  
                when "000111000010" => char <= "00100000";	--  
                when "000111000011" => char <= "00100000";	--  
                when "000111000100" => char <= "00100000";	--  
                when "000111000101" => char <= "01000000";	-- @
                when "000111000110" => char <= "01000000";	-- @
                when "000111000111" => char <= "01000000";	-- @
                when "000111001000" => char <= "01000000";	-- @
                when "000111001001" => char <= "01000000";	-- @
                when "000111001010" => char <= "01000000";	-- @
                when "000111001011" => char <= "01000000";	-- @
                when "000111001100" => char <= "01000000";	-- @
                when "000111001101" => char <= "01000000";	-- @
                when "000111001110" => char <= "01000000";	-- @

                when "001000000001" => char <= "00100000";	--  
                when "001000000010" => char <= "00100000";	--  
                when "001000000011" => char <= "00100000";	--  
                when "001000000100" => char <= "00100000";	--  
                when "001000000101" => char <= "00100000";	--  
                when "001000000110" => char <= "00100000";	--  
                when "001000000111" => char <= "01000000";	-- @
                when "001000001000" => char <= "01000000";	-- @
                when "001000001001" => char <= "01000000";	-- @
                when "001000001010" => char <= "01000000";	-- @
                when "001000001011" => char <= "01000000";	-- @
                when "001000001100" => char <= "01000000";	-- @

                when "001001000001" => char <= "00100000";	--  
                when "001001000010" => char <= "00100000";	--  
                when "001001000011" => char <= "00100000";	--  
                when "001001000100" => char <= "00100000";	--  
                when "001001000101" => char <= "00100000";	--  
                when "001001000110" => char <= "00100000";	--  
                when "001001000111" => char <= "00100000";	--  
                when "001001001000" => char <= "00100000";	--  
                when "001001001001" => char <= "01000000";	-- @
                when "001001001010" => char <= "01000000";	-- @

                when         others => char <= "00000000";
            end case;
        end if;
    end process;

end;
