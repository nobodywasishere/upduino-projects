library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity text_buffer is
	port(
        clk : in std_logic;
        row : in unsigned(5 downto 0);
        col : in unsigned(5 downto 0);
        char : out unsigned(7 downto 0)
	);
end text_buffer;

architecture synth of text_buffer is

    signal addr : unsigned (11 downto 0) := (others => '0');

begin

    addr <= row & col;

    process (clk) begin
        if (rising_edge(clk)) then
            case addr is

                when "000000000000" => char <= "01000001"; -- A
                when "000000000001" => char <= "01000010"; -- B
                when "000000000010" => char <= "01000011"; -- C
                when "000000000011" => char <= "01000100"; -- D
                when "000000000100" => char <= "01000101"; -- E
                when "000000000101" => char <= "01000110"; -- F
                when "000000000110" => char <= "01000111"; -- G
                when "000000000111" => char <= "01001000"; -- H
                when "000000001000" => char <= "01001001"; -- I
                when "000000001001" => char <= "01001010"; -- J
                when "000000001010" => char <= "01001011"; -- K
                when "000000001011" => char <= "01001100"; -- L
                when "000000001100" => char <= "01001101"; -- M
                when "000000001101" => char <= "01001110"; -- N
                when "000000001110" => char <= "01001111"; -- O
                when "000000001111" => char <= "01010000"; -- P
                when "000000010000" => char <= "01010001"; -- Q
                when "000000010001" => char <= "01010010"; -- R
                when "000000010010" => char <= "01010011"; -- S
                when "000000010011" => char <= "01010100"; -- T
                when "000000010100" => char <= "01010101"; -- U
                when "000000010101" => char <= "01010110"; -- V
                when "000000010110" => char <= "01010111"; -- W
                when "000000010111" => char <= "01011000"; -- X
                when "000000011000" => char <= "01011001"; -- Y
                when "000000011001" => char <= "01011010"; -- Z
                when "000000011010" => char <= "01011011"; --
                when "000000011011" => char <= "01011100"; --
                when "000000011100" => char <= "01011101"; --
                when "000000011101" => char <= "01011110"; --
                when "000000011110" => char <= "01011111"; --
                when "000000011111" => char <= "01011111"; --
                when "000000100000" => char <= "00000000";
                when "000000100001" => char <= "00000000";
                when "000000100010" => char <= "00000000";
                when "000000100011" => char <= "00000000";
                when "000000100100" => char <= "00000000";
                when "000000100101" => char <= "00000000";
                when "000000100110" => char <= "00000000";
                when "000000100111" => char <= "00000000";
                when "000000101000" => char <= "00000000";

                -- when "000001000000" => char <= "00000000";
                -- when "000001000001" => char <= "00000000";
                -- when "000001000010" => char <= "00000000";
                -- when "000001000011" => char <= "00000000";
                -- when "000001000100" => char <= "00000000";
                -- when "000001000101" => char <= "00000000";
                -- when "000001000110" => char <= "00000000";
                -- when "000001000111" => char <= "00000000";
                -- when "000001001000" => char <= "00000000";
                -- when "000001001001" => char <= "00000000";
                -- when "000001001010" => char <= "00000000";
                -- when "000001001011" => char <= "00000000";
                -- when "000001001100" => char <= "00000000";
                -- when "000001001101" => char <= "00000000";
                -- when "000001001110" => char <= "00000000";
                -- when "000001001111" => char <= "00000000";
                -- when "000001010000" => char <= "00000000";
                -- when "000001010001" => char <= "00000000";
                -- when "000001010010" => char <= "00000000";
                -- when "000001010011" => char <= "00000000";
                -- when "000001010100" => char <= "00000000";
                -- when "000001010101" => char <= "00000000";
                -- when "000001010110" => char <= "00000000";
                -- when "000001010111" => char <= "00000000";
                -- when "000001011000" => char <= "00000000";
                -- when "000001011001" => char <= "00000000";
                -- when "000001011010" => char <= "00000000";
                -- when "000001011011" => char <= "00000000";
                -- when "000001011100" => char <= "00000000";
                -- when "000001011101" => char <= "00000000";
                -- when "000001011110" => char <= "00000000";
                -- when "000001011111" => char <= "00000000";
                -- when "000001100000" => char <= "00000000";
                -- when "000001100001" => char <= "00000000";
                -- when "000001100010" => char <= "00000000";
                -- when "000001100011" => char <= "00000000";
                -- when "000001100100" => char <= "00000000";
                -- when "000001100101" => char <= "00000000";
                -- when "000001100110" => char <= "00000000";
                -- when "000001100111" => char <= "00000000";
                -- when "000001101000" => char <= "00000000";

                when "000010000000" => char <= "01000001";
                when "000010000001" => char <= "01000011";
                when "000010000010" => char <= "01000011";
                when "000010000011" => char <= "01001111";
                when "000010000100" => char <= "01010010";
                when "000010000101" => char <= "01000100";
                when "000010000110" => char <= "01001001";
                when "000010000111" => char <= "01001110";
                when "000010001000" => char <= "01000111";
                when "000010001001" => char <= "00000000";
                when "000010001010" => char <= "01010100";
                when "000010001011" => char <= "01001111";
                when "000010001100" => char <= "00000000";
                when "000010001101" => char <= "01000001";
                when "000010001110" => char <= "01001100";
                when "000010001111" => char <= "01001100";
                when "000010010000" => char <= "00000000";
                when "000010010001" => char <= "01001011";
                when "000010010010" => char <= "01001110";
                when "000010010011" => char <= "01001111";
                when "000010010100" => char <= "01010111";
                when "000010010101" => char <= "01001110";
                when "000010010110" => char <= "00000000";
                when "000010010111" => char <= "01001100";
                when "000010011000" => char <= "01000001";
                when "000010011001" => char <= "01010111";
                when "000010011010" => char <= "01010011";
                when "000010011011" => char <= "00000000";
                when "000010011100" => char <= "01001111";
                when "000010011101" => char <= "01000110";
                when "000010011110" => char <= "00000000";
                when "000010011111" => char <= "01000001";
                when "000010100000" => char <= "01010110";
                when "000010100001" => char <= "01001001";
                when "000010100010" => char <= "01000001";
                when "000010100011" => char <= "01010100";
                when "000010100100" => char <= "01001001";
                when "000010100101" => char <= "01001111";
                when "000010100110" => char <= "01001110";
                when "000010100111" => char <= "00000000";
                when "000010101000" => char <= "00000000";

                when "000011000000" => char <= "01010100";
                when "000011000001" => char <= "01001000";
                when "000011000010" => char <= "01000101";
                when "000011000011" => char <= "01010010";
                when "000011000100" => char <= "01000101";
                when "000011000101" => char <= "00000000";
                when "000011000110" => char <= "01001001";
                when "000011000111" => char <= "01010011";
                when "000011001000" => char <= "00000000";
                when "000011001001" => char <= "01001110";
                when "000011001010" => char <= "01001111";
                when "000011001011" => char <= "00000000";
                when "000011001100" => char <= "01010111";
                when "000011001101" => char <= "01000001";
                when "000011001110" => char <= "01011001";
                when "000011001111" => char <= "00000000";
                when "000011010000" => char <= "01010100";
                when "000011010001" => char <= "01001000";
                when "000011010010" => char <= "01000001";
                when "000011010011" => char <= "01010100";
                when "000011010100" => char <= "00000000";
                when "000011010101" => char <= "01000001";
                when "000011010110" => char <= "00000000";
                when "000011010111" => char <= "01000010";
                when "000011011000" => char <= "01000101";
                when "000011011001" => char <= "01000101";
                when "000011011010" => char <= "00000000";
                when "000011011011" => char <= "01010011";
                when "000011011100" => char <= "01001000";
                when "000011011101" => char <= "01001111";
                when "000011011110" => char <= "01010101";
                when "000011011111" => char <= "01001100";
                when "000011100000" => char <= "01000100";
                when "000011100001" => char <= "00000000";
                when "000011100010" => char <= "01000010";
                when "000011100011" => char <= "01000101";
                when "000011100100" => char <= "00000000";
                when "000011100101" => char <= "00000000";
                when "000011100110" => char <= "00000000";
                when "000011100111" => char <= "00000000";
                when "000011101000" => char <= "00000000";

                when "000100000000" => char <= "01000001";
                when "000100000001" => char <= "01000010";
                when "000100000010" => char <= "01001100";
                when "000100000011" => char <= "01000101";
                when "000100000100" => char <= "00000000";
                when "000100000101" => char <= "01010100";
                when "000100000110" => char <= "01001111";
                when "000100000111" => char <= "00000000";
                when "000100001000" => char <= "01000110";
                when "000100001001" => char <= "01001100";
                when "000100001010" => char <= "01011001";
                when "000100001011" => char <= "00000000";
                when "000100001100" => char <= "00000000";
                when "000100001101" => char <= "00000000";
                when "000100001110" => char <= "00000000";
                when "000100001111" => char <= "00000000";
                when "000100010000" => char <= "00000000";
                when "000100010001" => char <= "00000000";
                when "000100010010" => char <= "00000000";
                when "000100010011" => char <= "00000000";
                when "000100010100" => char <= "00000000";
                when "000100010101" => char <= "00000000";
                when "000100010110" => char <= "00000000";
                when "000100010111" => char <= "00000000";
                when "000100011000" => char <= "00000000";
                when "000100011001" => char <= "00000000";
                when "000100011010" => char <= "00000000";
                when "000100011011" => char <= "00000000";
                when "000100011100" => char <= "00000000";
                when "000100011101" => char <= "00000000";
                when "000100011110" => char <= "00000000";
                when "000100011111" => char <= "00000000";
                when "000100100000" => char <= "00000000";
                when "000100100001" => char <= "00000000";
                when "000100100010" => char <= "00000000";
                when "000100100011" => char <= "00000000";
                when "000100100100" => char <= "00000000";
                when "000100100101" => char <= "00000000";
                when "000100100110" => char <= "00000000";
                when "000100100111" => char <= "00000000";
                when "000100101000" => char <= "00000000";

                -- when "000101000000" => char <= "00000000";
                -- when "000101000001" => char <= "00000000";
                -- when "000101000010" => char <= "00000000";
                -- when "000101000011" => char <= "00000000";
                -- when "000101000100" => char <= "00000000";
                -- when "000101000101" => char <= "00000000";
                -- when "000101000110" => char <= "00000000";
                -- when "000101000111" => char <= "00000000";
                -- when "000101001000" => char <= "00000000";
                -- when "000101001001" => char <= "00000000";
                -- when "000101001010" => char <= "00000000";
                -- when "000101001011" => char <= "00000000";
                -- when "000101001100" => char <= "00000000";
                -- when "000101001101" => char <= "00000000";
                -- when "000101001110" => char <= "00000000";
                -- when "000101001111" => char <= "00000000";
                -- when "000101010000" => char <= "00000000";
                -- when "000101010001" => char <= "00000000";
                -- when "000101010010" => char <= "00000000";
                -- when "000101010011" => char <= "00000000";
                -- when "000101010100" => char <= "00000000";
                -- when "000101010101" => char <= "00000000";
                -- when "000101010110" => char <= "00000000";
                -- when "000101010111" => char <= "00000000";
                -- when "000101011000" => char <= "00000000";
                -- when "000101011001" => char <= "00000000";
                -- when "000101011010" => char <= "00000000";
                -- when "000101011011" => char <= "00000000";
                -- when "000101011100" => char <= "00000000";
                -- when "000101011101" => char <= "00000000";
                -- when "000101011110" => char <= "00000000";
                -- when "000101011111" => char <= "00000000";
                -- when "000101100000" => char <= "00000000";
                -- when "000101100001" => char <= "00000000";
                -- when "000101100010" => char <= "00000000";
                -- when "000101100011" => char <= "00000000";
                -- when "000101100100" => char <= "00000000";
                -- when "000101100101" => char <= "00000000";
                -- when "000101100110" => char <= "00000000";
                -- when "000101100111" => char <= "00000000";
                -- when "000101101000" => char <= "00000000";

                when "000110000000" => char <= "01001001";
                when "000110000001" => char <= "01010100";
                when "000110000010" => char <= "01010011";
                when "000110000011" => char <= "00000000";
                when "000110000100" => char <= "01010111";
                when "000110000101" => char <= "01001001";
                when "000110000110" => char <= "01001110";
                when "000110000111" => char <= "01000111";
                when "000110001000" => char <= "01010011";
                when "000110001001" => char <= "00000000";
                when "000110001010" => char <= "01000001";
                when "000110001011" => char <= "01010010";
                when "000110001100" => char <= "01000101";
                when "000110001101" => char <= "00000000";
                when "000110001110" => char <= "01010100";
                when "000110001111" => char <= "01001111";
                when "000110010000" => char <= "01001111";
                when "000110010001" => char <= "00000000";
                when "000110010010" => char <= "01010011";
                when "000110010011" => char <= "01001101";
                when "000110010100" => char <= "01000001";
                when "000110010101" => char <= "01001100";
                when "000110010110" => char <= "01001100";
                when "000110010111" => char <= "00000000";
                when "000110011000" => char <= "01010100";
                when "000110011001" => char <= "01001111";
                when "000110011010" => char <= "00000000";
                when "000110011011" => char <= "01000111";
                when "000110011100" => char <= "01000101";
                when "000110011101" => char <= "01010100";
                when "000110011110" => char <= "00000000";
                when "000110011111" => char <= "01001001";
                when "000110100000" => char <= "01010100";
                when "000110100001" => char <= "01010011";
                when "000110100010" => char <= "00000000";
                when "000110100011" => char <= "00000000";
                when "000110100100" => char <= "00000000";
                when "000110100101" => char <= "00000000";
                when "000110100110" => char <= "00000000";
                when "000110100111" => char <= "00000000";
                when "000110101000" => char <= "00000000";

                when "000111000000" => char <= "01000110";
                when "000111000001" => char <= "01000001";
                when "000111000010" => char <= "01010100";
                when "000111000011" => char <= "00000000";
                when "000111000100" => char <= "01001100";
                when "000111000101" => char <= "01001001";
                when "000111000110" => char <= "01010100";
                when "000111000111" => char <= "01010100";
                when "000111001000" => char <= "01001100";
                when "000111001001" => char <= "01000101";
                when "000111001010" => char <= "00000000";
                when "000111001011" => char <= "01000010";
                when "000111001100" => char <= "01001111";
                when "000111001101" => char <= "01000100";
                when "000111001110" => char <= "01011001";
                when "000111001111" => char <= "00000000";
                when "000111010000" => char <= "01001111";
                when "000111010001" => char <= "01000110";
                when "000111010010" => char <= "01000110";
                when "000111010011" => char <= "00000000";
                when "000111010100" => char <= "01010100";
                when "000111010101" => char <= "01001000";
                when "000111010110" => char <= "01000101";
                when "000111010111" => char <= "00000000";
                when "000111011000" => char <= "01000111";
                when "000111011001" => char <= "01010010";
                when "000111011010" => char <= "01001111";
                when "000111011011" => char <= "01010101";
                when "000111011100" => char <= "01001110";
                when "000111011101" => char <= "01000100";
                when "000111011110" => char <= "00000000";
                when "000111011111" => char <= "00000000";
                when "000111100000" => char <= "00000000";
                when "000111100001" => char <= "00000000";
                when "000111100010" => char <= "00000000";
                when "000111100011" => char <= "00000000";
                when "000111100100" => char <= "00000000";
                when "000111100101" => char <= "00000000";
                when "000111100110" => char <= "00000000";
                when "000111100111" => char <= "00000000";
                when "000111101000" => char <= "00000000";

                -- when "001000000000" => char <= "00000000";
                -- when "001000000001" => char <= "00000000";
                -- when "001000000010" => char <= "00000000";
                -- when "001000000011" => char <= "00000000";
                -- when "001000000100" => char <= "00000000";
                -- when "001000000101" => char <= "00000000";
                -- when "001000000110" => char <= "00000000";
                -- when "001000000111" => char <= "00000000";
                -- when "001000001000" => char <= "00000000";
                -- when "001000001001" => char <= "00000000";
                -- when "001000001010" => char <= "00000000";
                -- when "001000001011" => char <= "00000000";
                -- when "001000001100" => char <= "00000000";
                -- when "001000001101" => char <= "00000000";
                -- when "001000001110" => char <= "00000000";
                -- when "001000001111" => char <= "00000000";
                -- when "001000010000" => char <= "00000000";
                -- when "001000010001" => char <= "00000000";
                -- when "001000010010" => char <= "00000000";
                -- when "001000010011" => char <= "00000000";
                -- when "001000010100" => char <= "00000000";
                -- when "001000010101" => char <= "00000000";
                -- when "001000010110" => char <= "00000000";
                -- when "001000010111" => char <= "00000000";
                -- when "001000011000" => char <= "00000000";
                -- when "001000011001" => char <= "00000000";
                -- when "001000011010" => char <= "00000000";
                -- when "001000011011" => char <= "00000000";
                -- when "001000011100" => char <= "00000000";
                -- when "001000011101" => char <= "00000000";
                -- when "001000011110" => char <= "00000000";
                -- when "001000011111" => char <= "00000000";
                -- when "001000100000" => char <= "00000000";
                -- when "001000100001" => char <= "00000000";
                -- when "001000100010" => char <= "00000000";
                -- when "001000100011" => char <= "00000000";
                -- when "001000100100" => char <= "00000000";
                -- when "001000100101" => char <= "00000000";
                -- when "001000100110" => char <= "00000000";
                -- when "001000100111" => char <= "00000000";
                -- when "001000101000" => char <= "00000000";
                --
                when "001001000000" => char <= "01010100";
                when "001001000001" => char <= "01001000";
                when "001001000010" => char <= "01000101";
                when "001001000011" => char <= "00000000";
                when "001001000100" => char <= "01000010";
                when "001001000101" => char <= "01000101";
                when "001001000110" => char <= "01000101";
                when "001001000111" => char <= "00000000";
                when "001001001000" => char <= "01001111";
                when "001001001001" => char <= "01000110";
                when "001001001010" => char <= "00000000";
                when "001001001011" => char <= "01000011";
                when "001001001100" => char <= "01001111";
                when "001001001101" => char <= "01010101";
                when "001001001110" => char <= "01010010";
                when "001001001111" => char <= "01010011";
                when "001001010000" => char <= "01000101";
                when "001001010001" => char <= "00000000";
                when "001001010010" => char <= "01000110";
                when "001001010011" => char <= "01001100";
                when "001001010100" => char <= "01001001";
                when "001001010101" => char <= "01000101";
                when "001001010110" => char <= "01010011";
                when "001001010111" => char <= "00000000";
                when "001001011000" => char <= "01000001";
                when "001001011001" => char <= "01001110";
                when "001001011010" => char <= "01011001";
                when "001001011011" => char <= "01010111";
                when "001001011100" => char <= "01000001";
                when "001001011101" => char <= "01011001";
                when "001001011110" => char <= "01010011";
                when "001001011111" => char <= "00000000";
                when "001001100000" => char <= "00000000";
                when "001001100001" => char <= "00000000";
                when "001001100010" => char <= "00000000";
                when "001001100011" => char <= "00000000";
                when "001001100100" => char <= "00000000";
                when "001001100101" => char <= "00000000";
                when "001001100110" => char <= "00000000";
                when "001001100111" => char <= "00000000";
                when "001001101000" => char <= "00000000";
                --
                when "001010000000" => char <= "01000010";
                when "001010000001" => char <= "01000101";
                when "001010000010" => char <= "01000011";
                when "001010000011" => char <= "01000001";
                when "001010000100" => char <= "01010101";
                when "001010000101" => char <= "01010011";
                when "001010000110" => char <= "01000101";
                when "001010000111" => char <= "00000000";
                when "001010001000" => char <= "01000010";
                when "001010001001" => char <= "01000101";
                when "001010001010" => char <= "01000101";
                when "001010001011" => char <= "01010011";
                when "001010001100" => char <= "00000000";
                when "001010001101" => char <= "01000100";
                when "001010001110" => char <= "01001111";
                when "001010001111" => char <= "01001110";
                when "001010010000" => char <= "01010100";
                when "001010010001" => char <= "00000000";
                when "001010010010" => char <= "01000011";
                when "001010010011" => char <= "01000001";
                when "001010010100" => char <= "01010010";
                when "001010010101" => char <= "01000101";
                when "001010010110" => char <= "00000000";
                when "001010010111" => char <= "01010111";
                when "001010011000" => char <= "01001000";
                when "001010011001" => char <= "01000001";
                when "001010011010" => char <= "01010100";
                when "001010011011" => char <= "00000000";
                when "001010011100" => char <= "01001000";
                when "001010011101" => char <= "01010101";
                when "001010011110" => char <= "01001101";
                when "001010011111" => char <= "01000001";
                when "001010100000" => char <= "01001110";
                when "001010100001" => char <= "01010011";
                when "001010100010" => char <= "00000000";
                when "001010100011" => char <= "00000000";
                when "001010100100" => char <= "00000000";
                when "001010100101" => char <= "00000000";
                when "001010100110" => char <= "00000000";
                when "001010100111" => char <= "00000000";
                when "001010101000" => char <= "00000000";
                --
                when "001011000000" => char <= "01010100";
                when "001011000001" => char <= "01001000";
                when "001011000010" => char <= "01001001";
                when "001011000011" => char <= "01001110";
                when "001011000100" => char <= "01001011";
                when "001011000101" => char <= "00000000";
                when "001011000110" => char <= "01001001";
                when "001011000111" => char <= "01010011";
                when "001011001000" => char <= "00000000";
                when "001011001001" => char <= "01001001";
                when "001011001010" => char <= "01001101";
                when "001011001011" => char <= "01010000";
                when "001011001100" => char <= "01001111";
                when "001011001101" => char <= "01010011";
                when "001011001110" => char <= "01010011";
                when "001011001111" => char <= "01001001";
                when "001011010000" => char <= "01000010";
                when "001011010001" => char <= "01001100";
                when "001011010010" => char <= "01000101";
                when "001011010011" => char <= "00000000";
                when "001011010100" => char <= "00000000";
                when "001011010101" => char <= "00000000";
                when "001011010110" => char <= "00000000";
                when "001011010111" => char <= "00000000";
                when "001011011000" => char <= "00000000";
                when "001011011001" => char <= "00000000";
                when "001011011010" => char <= "00000000";
                when "001011011011" => char <= "00000000";
                when "001011011100" => char <= "00000000";
                when "001011011101" => char <= "00000000";
                when "001011011110" => char <= "00000000";
                when "001011011111" => char <= "00000000";
                when "001011100000" => char <= "00000000";
                when "001011100001" => char <= "00000000";
                when "001011100010" => char <= "00000000";
                when "001011100011" => char <= "00000000";
                when "001011100100" => char <= "00000000";
                when "001011100101" => char <= "00000000";
                when "001011100110" => char <= "00000000";
                when "001011100111" => char <= "00000000";
                when "001011101000" => char <= "00000000";
                --
                -- when "001100000000" => char <= "01000001";
                -- when "001100000001" => char <= "01000010";
                -- when "001100000010" => char <= "01000011";
                -- when "001100000011" => char <= "01000100";
                -- when "001100000100" => char <= "01000101";
                -- when "001100000101" => char <= "01000110";
                -- when "001100000110" => char <= "01000111";
                -- when "001100000111" => char <= "01001000";
                -- when "001100001000" => char <= "01001001";
                -- when "001100001001" => char <= "01001010";
                -- when "001100001010" => char <= "01001011";
                -- when "001100001011" => char <= "01001100";
                -- when "001100001100" => char <= "01001101";
                -- when "001100001101" => char <= "01001110";
                -- when "001100001110" => char <= "01001111";
                -- when "001100001111" => char <= "01010000";
                -- when "001100010000" => char <= "01010001";
                -- when "001100010001" => char <= "01010010";
                -- when "001100010010" => char <= "01010011";
                -- when "001100010011" => char <= "01010100";
                -- when "001100010100" => char <= "01010101";
                -- when "001100010101" => char <= "01010110";
                -- when "001100010110" => char <= "01010111";
                -- when "001100010111" => char <= "01011000";
                -- when "001100011000" => char <= "01011001";
                -- when "001100011001" => char <= "01011010";
                -- when "001100011010" => char <= "01011011";
                -- when "001100011011" => char <= "01011100";
                -- when "001100011100" => char <= "01011101";
                -- when "001100011101" => char <= "01011110";
                -- when "001100011110" => char <= "01011111";
                -- when "001100011111" => char <= "01011111";
                -- when "001100100000" => char <= "00000000";
                -- when "001100100001" => char <= "00000000";
                -- when "001100100010" => char <= "00000000";
                -- when "001100100011" => char <= "00000000";
                -- when "001100100100" => char <= "00000000";
                -- when "001100100101" => char <= "00000000";
                -- when "001100100110" => char <= "00000000";
                -- when "001100100111" => char <= "00000000";
                -- when "001100101000" => char <= "00000000";
                --
                -- when "001101000000" => char <= "01000001";
                -- when "001101000001" => char <= "01000010";
                -- when "001101000010" => char <= "01000011";
                -- when "001101000011" => char <= "01000100";
                -- when "001101000100" => char <= "01000101";
                -- when "001101000101" => char <= "01000110";
                -- when "001101000110" => char <= "01000111";
                -- when "001101000111" => char <= "01001000";
                -- when "001101001000" => char <= "01001001";
                -- when "001101001001" => char <= "01001010";
                -- when "001101001010" => char <= "01001011";
                -- when "001101001011" => char <= "01001100";
                -- when "001101001100" => char <= "01001101";
                -- when "001101001101" => char <= "01001110";
                -- when "001101001110" => char <= "01001111";
                -- when "001101001111" => char <= "01010000";
                -- when "001101010000" => char <= "01010001";
                -- when "001101010001" => char <= "01010010";
                -- when "001101010010" => char <= "01010011";
                -- when "001101010011" => char <= "01010100";
                -- when "001101010100" => char <= "01010101";
                -- when "001101010101" => char <= "01010110";
                -- when "001101010110" => char <= "01010111";
                -- when "001101010111" => char <= "01011000";
                -- when "001101011000" => char <= "01011001";
                -- when "001101011001" => char <= "01011010";
                -- when "001101011010" => char <= "01011011";
                -- when "001101011011" => char <= "01011100";
                -- when "001101011100" => char <= "01011101";
                -- when "001101011101" => char <= "01011110";
                -- when "001101011110" => char <= "01011111";
                -- when "001101011111" => char <= "01011111";
                -- when "001101100000" => char <= "00000000";
                -- when "001101100001" => char <= "00000000";
                -- when "001101100010" => char <= "00000000";
                -- when "001101100011" => char <= "00000000";
                -- when "001101100100" => char <= "00000000";
                -- when "001101100101" => char <= "00000000";
                -- when "001101100110" => char <= "00000000";
                -- when "001101100111" => char <= "00000000";
                -- when "001101101000" => char <= "00000000";
                --
                -- when "001110000000" => char <= "01000001";
                -- when "001110000001" => char <= "01000010";
                -- when "001110000010" => char <= "01000011";
                -- when "001110000011" => char <= "01000100";
                -- when "001110000100" => char <= "01000101";
                -- when "001110000101" => char <= "01000110";
                -- when "001110000110" => char <= "01000111";
                -- when "001110000111" => char <= "01001000";
                -- when "001110001000" => char <= "01001001";
                -- when "001110001001" => char <= "01001010";
                -- when "001110001010" => char <= "01001011";
                -- when "001110001011" => char <= "01001100";
                -- when "001110001100" => char <= "01001101";
                -- when "001110001101" => char <= "01001110";
                -- when "001110001110" => char <= "01001111";
                -- when "001110001111" => char <= "01010000";
                -- when "001110010000" => char <= "01010001";
                -- when "001110010001" => char <= "01010010";
                -- when "001110010010" => char <= "01010011";
                -- when "001110010011" => char <= "01010100";
                -- when "001110010100" => char <= "01010101";
                -- when "001110010101" => char <= "01010110";
                -- when "001110010110" => char <= "01010111";
                -- when "001110010111" => char <= "01011000";
                -- when "001110011000" => char <= "01011001";
                -- when "001110011001" => char <= "01011010";
                -- when "001110011010" => char <= "01011011";
                -- when "001110011011" => char <= "01011100";
                -- when "001110011100" => char <= "01011101";
                -- when "001110011101" => char <= "01011110";
                -- when "001110011110" => char <= "01011111";
                -- when "001110011111" => char <= "01011111";
                -- when "001110100000" => char <= "00000000";
                -- when "001110100001" => char <= "00000000";
                -- when "001110100010" => char <= "00000000";
                -- when "001110100011" => char <= "00000000";
                -- when "001110100100" => char <= "00000000";
                -- when "001110100101" => char <= "00000000";
                -- when "001110100110" => char <= "00000000";
                -- when "001110100111" => char <= "00000000";
                -- when "001110101000" => char <= "00000000";
                --
                -- when "001111000000" => char <= "01000001";
                -- when "001111000001" => char <= "01000010";
                -- when "001111000010" => char <= "01000011";
                -- when "001111000011" => char <= "01000100";
                -- when "001111000100" => char <= "01000101";
                -- when "001111000101" => char <= "01000110";
                -- when "001111000110" => char <= "01000111";
                -- when "001111000111" => char <= "01001000";
                -- when "001111001000" => char <= "01001001";
                -- when "001111001001" => char <= "01001010";
                -- when "001111001010" => char <= "01001011";
                -- when "001111001011" => char <= "01001100";
                -- when "001111001100" => char <= "01001101";
                -- when "001111001101" => char <= "01001110";
                -- when "001111001110" => char <= "01001111";
                -- when "001111001111" => char <= "01010000";
                -- when "001111010000" => char <= "01010001";
                -- when "001111010001" => char <= "01010010";
                -- when "001111010010" => char <= "01010011";
                -- when "001111010011" => char <= "01010100";
                -- when "001111010100" => char <= "01010101";
                -- when "001111010101" => char <= "01010110";
                -- when "001111010110" => char <= "01010111";
                -- when "001111010111" => char <= "01011000";
                -- when "001111011000" => char <= "01011001";
                -- when "001111011001" => char <= "01011010";
                -- when "001111011010" => char <= "01011011";
                -- when "001111011011" => char <= "01011100";
                -- when "001111011100" => char <= "01011101";
                -- when "001111011101" => char <= "01011110";
                -- when "001111011110" => char <= "01011111";
                -- when "001111011111" => char <= "01011111";
                -- when "001111100000" => char <= "00000000";
                -- when "001111100001" => char <= "00000000";
                -- when "001111100010" => char <= "00000000";
                -- when "001111100011" => char <= "00000000";
                -- when "001111100100" => char <= "00000000";
                -- when "001111100101" => char <= "00000000";
                -- when "001111100110" => char <= "00000000";
                -- when "001111100111" => char <= "00000000";
                -- when "001111101000" => char <= "00000000";

                when         others => char <= "00000000";
            end case;
        end if;
    end process;

end;
