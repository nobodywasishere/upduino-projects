library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;


entity text_font is
	port(
        clk : in std_logic;
        char : in unsigned(7 downto 0);
        row : in unsigned(2 downto 0);
        col : in unsigned(2 downto 0);
        lum : out std_logic
	);
end text_font;

architecture synth of text_font is

    signal addr : unsigned(10 downto 0) := (others => '0');
    signal mem : unsigned(7 downto 0);

begin

    addr <= char & row;
    lum <= mem(to_integer(col));

    process (clk) begin
        if (rising_edge(clk)) then
            case addr is

                -- A  01000001
                when "01000001000" => mem <= "00011000";
                when "01000001001" => mem <= "00111100";
                when "01000001010" => mem <= "01100110";
                when "01000001011" => mem <= "01111110";
                when "01000001100" => mem <= "01100110";
                when "01000001101" => mem <= "01100110";
                when "01000001110" => mem <= "01100110";
                when "01000001111" => mem <= "00000000";

                -- B  01000010
                when "01000010000" => mem <= "00111110";
                when "01000010001" => mem <= "01100110";
                when "01000010010" => mem <= "01100110";
                when "01000010011" => mem <= "00111110";
                when "01000010100" => mem <= "01100110";
                when "01000010101" => mem <= "01100110";
                when "01000010110" => mem <= "00111110";
                when "01000010111" => mem <= "00000000";

                -- C  01000011
                when "01000011000" => mem <= "00111100";
                when "01000011001" => mem <= "01100110";
                when "01000011010" => mem <= "00000110";
                when "01000011011" => mem <= "00000110";
                when "01000011100" => mem <= "00000110";
                when "01000011101" => mem <= "01100110";
                when "01000011110" => mem <= "00111100";
                when "01000011111" => mem <= "00000000";

                -- D  01000100
                when "01000100000" => mem <= "00011110";
                when "01000100001" => mem <= "00110110";
                when "01000100010" => mem <= "01100110";
                when "01000100011" => mem <= "01100110";
                when "01000100100" => mem <= "01100110";
                when "01000100101" => mem <= "00110110";
                when "01000100110" => mem <= "00011110";
                when "01000100111" => mem <= "00000000";

                -- E  01000101
                when "01000101000" => mem <= "01111110";
                when "01000101001" => mem <= "00000110";
                when "01000101010" => mem <= "00000110";
                when "01000101011" => mem <= "00011110";
                when "01000101100" => mem <= "00000110";
                when "01000101101" => mem <= "00000110";
                when "01000101110" => mem <= "01111110";
                when "01000101111" => mem <= "00000000";

                -- F  01000110
                when "01000110000" => mem <= "01111110";
                when "01000110001" => mem <= "00000110";
                when "01000110010" => mem <= "00000110";
                when "01000110011" => mem <= "00011110";
                when "01000110100" => mem <= "00000110";
                when "01000110101" => mem <= "00000110";
                when "01000110110" => mem <= "00000110";
                when "01000110111" => mem <= "00000000";

                -- G  01000111
                when "01000111000" => mem <= "00111100";
                when "01000111001" => mem <= "01100110";
                when "01000111010" => mem <= "00000110";
                when "01000111011" => mem <= "01110110";
                when "01000111100" => mem <= "01100110";
                when "01000111101" => mem <= "01100110";
                when "01000111110" => mem <= "00111100";
                when "01000111111" => mem <= "00000000";

                -- H  01001000
                when "01001000000" => mem <= "01100110";
                when "01001000001" => mem <= "01100110";
                when "01001000010" => mem <= "01100110";
                when "01001000011" => mem <= "01111110";
                when "01001000100" => mem <= "01100110";
                when "01001000101" => mem <= "01100110";
                when "01001000110" => mem <= "01100110";
                when "01001000111" => mem <= "00000000";

                -- I  01001001
                when "01001001000" => mem <= "00111100";
                when "01001001001" => mem <= "00011000";
                when "01001001010" => mem <= "00011000";
                when "01001001011" => mem <= "00011000";
                when "01001001100" => mem <= "00011000";
                when "01001001101" => mem <= "00011000";
                when "01001001110" => mem <= "00111100";
                when "01001001111" => mem <= "00000000";

                -- J  01001010
                when "01001010000" => mem <= "01111000";
                when "01001010001" => mem <= "00110000";
                when "01001010010" => mem <= "00110000";
                when "01001010011" => mem <= "00110000";
                when "01001010100" => mem <= "00110000";
                when "01001010101" => mem <= "00110110";
                when "01001010110" => mem <= "00011100";
                when "01001010111" => mem <= "00000000";

                -- K  01001011
                when "01001011000" => mem <= "01100110";
                when "01001011001" => mem <= "00110110";
                when "01001011010" => mem <= "00011110";
                when "01001011011" => mem <= "00001110";
                when "01001011100" => mem <= "00011110";
                when "01001011101" => mem <= "00110110";
                when "01001011110" => mem <= "01100110";
                when "01001011111" => mem <= "00000000";

                -- L  01001100
                when "01001100000" => mem <= "00000110";
                when "01001100001" => mem <= "00000110";
                when "01001100010" => mem <= "00000110";
                when "01001100011" => mem <= "00000110";
                when "01001100100" => mem <= "00000110";
                when "01001100101" => mem <= "00000110";
                when "01001100110" => mem <= "01111110";
                when "01001100111" => mem <= "00000000";

                -- M  01001101
                when "01001101000" => mem <= "01000110";
                when "01001101001" => mem <= "01101110";
                when "01001101010" => mem <= "01111110";
                when "01001101011" => mem <= "01010110";
                when "01001101100" => mem <= "01000110";
                when "01001101101" => mem <= "01000110";
                when "01001101110" => mem <= "01000110";
                when "01001101111" => mem <= "00000000";

                -- N  01001110
                when "01001110000" => mem <= "01100110";
                when "01001110001" => mem <= "01101110";
                when "01001110010" => mem <= "01111110";
                when "01001110011" => mem <= "01111110";
                when "01001110100" => mem <= "01110110";
                when "01001110101" => mem <= "01100110";
                when "01001110110" => mem <= "01100110";
                when "01001110111" => mem <= "00000000";

                -- O  01001111
                when "01001111000" => mem <= "00111100";
                when "01001111001" => mem <= "01100110";
                when "01001111010" => mem <= "01100110";
                when "01001111011" => mem <= "01100110";
                when "01001111100" => mem <= "01100110";
                when "01001111101" => mem <= "01100110";
                when "01001111110" => mem <= "00111100";
                when "01001111111" => mem <= "00000000";

                -- P  01010000
                when "01010000000" => mem <= "00111110";
                when "01010000001" => mem <= "01100110";
                when "01010000010" => mem <= "01100110";
                when "01010000011" => mem <= "00111110";
                when "01010000100" => mem <= "00000110";
                when "01010000101" => mem <= "00000110";
                when "01010000110" => mem <= "00000110";
                when "01010000111" => mem <= "00000000";

                -- Q  01010001
                when "01010001000" => mem <= "00111110";
                when "01010001001" => mem <= "01100110";
                when "01010001010" => mem <= "01100110";
                when "01010001011" => mem <= "01100110";
                when "01010001100" => mem <= "01100110";
                when "01010001101" => mem <= "00111100";
                when "01010001110" => mem <= "01110000";
                when "01010001111" => mem <= "00000000";

                -- R  01010010
                when "01010010000" => mem <= "00111110";
                when "01010010001" => mem <= "01100110";
                when "01010010010" => mem <= "01100110";
                when "01010010011" => mem <= "00111110";
                when "01010010100" => mem <= "00011110";
                when "01010010101" => mem <= "00110110";
                when "01010010110" => mem <= "01100110";
                when "01010010111" => mem <= "00000000";

                -- S  01010011
                when "01010011000" => mem <= "00111100";
                when "01010011001" => mem <= "01100110";
                when "01010011010" => mem <= "00000110";
                when "01010011011" => mem <= "00111100";
                when "01010011100" => mem <= "01100000";
                when "01010011101" => mem <= "01100110";
                when "01010011110" => mem <= "00111100";
                when "01010011111" => mem <= "00000000";

                -- T  01010100
                when "01010100000" => mem <= "01111110";
                when "01010100001" => mem <= "00011000";
                when "01010100010" => mem <= "00011000";
                when "01010100011" => mem <= "00011000";
                when "01010100100" => mem <= "00011000";
                when "01010100101" => mem <= "00011000";
                when "01010100110" => mem <= "00011000";
                when "01010100111" => mem <= "00000000";

                -- U  01010101
                when "01010101000" => mem <= "01100110";
                when "01010101001" => mem <= "01100110";
                when "01010101010" => mem <= "01100110";
                when "01010101011" => mem <= "01100110";
                when "01010101100" => mem <= "01100110";
                when "01010101101" => mem <= "01100110";
                when "01010101110" => mem <= "00111100";
                when "01010101111" => mem <= "00000000";

                -- V  01010110
                when "01010110000" => mem <= "01100110";
                when "01010110001" => mem <= "01100110";
                when "01010110010" => mem <= "01100110";
                when "01010110011" => mem <= "01100110";
                when "01010110100" => mem <= "01100110";
                when "01010110101" => mem <= "00111100";
                when "01010110110" => mem <= "00011000";
                when "01010110111" => mem <= "00000000";

                -- W  01010111
                when "01010111000" => mem <= "01000110";
                when "01010111001" => mem <= "01000110";
                when "01010111010" => mem <= "01000110";
                when "01010111011" => mem <= "01010110";
                when "01010111100" => mem <= "01111110";
                when "01010111101" => mem <= "01101110";
                when "01010111110" => mem <= "01000110";
                when "01010111111" => mem <= "00000000";

                -- X  01011000
                when "01011000000" => mem <= "01100110";
                when "01011000001" => mem <= "01100110";
                when "01011000010" => mem <= "00111100";
                when "01011000011" => mem <= "00011000";
                when "01011000100" => mem <= "00111100";
                when "01011000101" => mem <= "01100110";
                when "01011000110" => mem <= "01100110";
                when "01011000111" => mem <= "00000000";

                -- Y  01011001
                when "01011001000" => mem <= "01100110";
                when "01011001001" => mem <= "01100110";
                when "01011001010" => mem <= "01100110";
                when "01011001011" => mem <= "00111100";
                when "01011001100" => mem <= "00011000";
                when "01011001101" => mem <= "00011000";
                when "01011001110" => mem <= "00011000";
                when "01011001111" => mem <= "00000000";

                -- Z  01011010
                when "01011010000" => mem <= "01111110";
                when "01011010001" => mem <= "01100000";
                when "01011010010" => mem <= "00110000";
                when "01011010011" => mem <= "00011000";
                when "01011010100" => mem <= "00001100";
                when "01011010101" => mem <= "00000110";
                when "01011010110" => mem <= "01111110";
                when "01011010111" => mem <= "00000000";

                when        others => mem <= "00000000";
            end case;
        end if;
    end process;

end;
